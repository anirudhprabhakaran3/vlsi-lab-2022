*nmos characteristics
*


m0 drain0 gate 0 0 nfet1 w=6.4u l=1.8u ad=6.84p pd=10.8u as=6.84p ps=10.8u
m1 drain1 gate 0 0 nfet2 w=6.4u l=1.8u ad=6.84p pd=10.8u as=6.84p ps=10.8u
m2 drain2 gate 0 0 nfet3 w=6.4u l=1.8u ad=6.84p pd=10.8u as=6.84p ps=10.8u
m4 drain3 gate 0 0 nfet4 w=6.4u l=1.8u
R0 dd drain0 0.0001
R1 dd drain1 0.0001
R2 dd drain2 0.0001
R3 dd drain3 0.0001


*
.MODEL nfet1 NMOS LEVEL=1 LAMBDA=0.5
.MODEL nfet2 NMOS LEVEL=1 LAMBDA=1.0
.MODEL nfet3 NMOS LEVEL=1 LAMBDA=1.5
.MODEL nfet4 NMOS LEVEL=1 LAMBDA=0.0
*

* supply voltages
Vdd dd 0 dc 5
Vgg gate 0 dc 5


*
* analysis request
.dc vdd 0 10 0.1 vgg 0 5 1
.control
run
setplot dc1
plot (v(dd)-v(drain0))/0.0001
plot (v(dd)-v(drain1))/0.0001
plot (v(dd)-v(drain2))/0.0001
plot (v(dd)-v(drain3))/0.0001
*plot (v(dd)-v(drain0))/0.0001 (v(dd)-v(drain1))/0.0001 (v(dd)-v(drain2))/0.0001
.endc

.end

