magic
tech scmos
timestamp 1666709236
<< pwell >>
rect 0 29 28 32
rect 0 8 32 29
rect 18 6 32 8
<< nwell >>
rect 0 50 32 64
rect 0 32 28 50
<< polysilicon >>
rect 5 60 7 62
rect 23 60 25 62
rect 5 23 7 44
rect 23 23 25 44
rect 5 12 7 15
rect 23 12 25 15
<< ndiffusion >>
rect 0 21 5 23
rect 4 17 5 21
rect 0 15 5 17
rect 7 21 23 23
rect 7 17 13 21
rect 17 17 23 21
rect 7 15 23 17
rect 25 21 32 23
rect 25 17 28 21
rect 25 15 32 17
<< pdiffusion >>
rect 0 53 5 60
rect 4 49 5 53
rect 0 44 5 49
rect 7 44 23 60
rect 25 54 32 60
rect 25 44 28 54
<< metal1 >>
rect 0 64 32 72
rect 0 53 4 64
rect 28 30 32 50
rect 13 26 32 30
rect 13 21 17 26
rect 0 8 4 17
rect 28 8 32 17
rect 0 0 32 8
<< ntransistor >>
rect 5 15 7 23
rect 23 15 25 23
<< ptransistor >>
rect 5 44 7 60
rect 23 44 25 60
<< polycontact >>
rect 1 37 5 41
rect 19 37 23 41
<< ndcontact >>
rect 0 17 4 21
rect 13 17 17 21
rect 28 17 32 21
<< pdcontact >>
rect 0 49 4 53
rect 28 50 32 54
<< labels >>
rlabel metal1 15 68 15 68 5 vdd
rlabel polycontact 3 39 3 39 3 a
rlabel polycontact 21 39 21 39 1 b
rlabel metal1 15 3 15 3 1 vss
rlabel metal1 30 28 30 28 7 output
<< end >>
