magic
tech scmos
timestamp 1666019148
<< ab >>
rect -139 31 -75 77
rect 5 57 29 77
rect 7 53 29 57
rect -36 37 -30 39
rect -70 31 0 37
rect -139 27 0 31
rect -139 5 -75 27
rect -70 1 0 27
rect 5 5 29 53
rect -70 0 1 1
<< nwell >>
rect -141 60 -70 82
rect 0 60 34 82
rect -141 37 34 60
<< pwell >>
rect -141 5 34 37
rect -92 0 34 5
<< poly >>
rect -129 67 -118 69
rect -129 65 -127 67
rect -133 63 -127 65
rect -120 64 -118 67
rect -133 61 -131 63
rect -129 61 -127 63
rect -133 59 -127 61
rect -100 63 -94 65
rect -86 64 -84 69
rect -100 61 -98 63
rect -96 61 -94 63
rect -106 56 -104 61
rect -100 59 -94 61
rect -96 56 -94 59
rect 14 62 20 64
rect 14 60 16 62
rect 18 60 20 62
rect 14 58 20 60
rect 14 55 16 58
rect -120 40 -118 43
rect -106 40 -104 43
rect -126 38 -118 40
rect -114 38 -104 40
rect -126 31 -124 38
rect -114 36 -112 38
rect -110 36 -108 38
rect -114 34 -108 36
rect -113 25 -111 34
rect -96 30 -94 43
rect -86 40 -84 43
rect -90 38 -84 40
rect -90 36 -88 38
rect -86 36 -84 38
rect -90 34 -84 36
rect -103 25 -101 30
rect -96 28 -91 30
rect -93 25 -91 28
rect -86 25 -84 34
rect 14 31 16 43
rect -126 10 -124 24
rect -113 14 -111 18
rect -103 10 -101 18
rect 14 20 16 25
rect -93 11 -91 16
rect -86 11 -84 16
rect -126 8 -101 10
<< ndif >>
rect -133 29 -126 31
rect -133 27 -131 29
rect -129 27 -126 29
rect -133 24 -126 27
rect -124 25 -115 31
rect 7 29 14 31
rect 7 27 9 29
rect 11 27 14 29
rect 7 25 14 27
rect 16 29 23 31
rect 16 27 19 29
rect 21 27 23 29
rect 16 25 23 27
rect -124 24 -113 25
rect -122 22 -113 24
rect -122 20 -120 22
rect -118 20 -113 22
rect -122 18 -113 20
rect -111 22 -103 25
rect -111 20 -108 22
rect -106 20 -103 22
rect -111 18 -103 20
rect -101 22 -93 25
rect -101 20 -98 22
rect -96 20 -93 22
rect -101 18 -93 20
rect -98 16 -93 18
rect -91 16 -86 25
rect -84 20 -77 25
rect -84 18 -81 20
rect -79 18 -77 20
rect -84 16 -77 18
<< pdif >>
rect 7 72 13 74
rect 7 70 9 72
rect 11 70 13 72
rect -125 49 -120 64
rect -127 47 -120 49
rect -127 45 -125 47
rect -123 45 -120 47
rect -127 43 -120 45
rect -118 62 -108 64
rect -118 60 -115 62
rect -113 60 -108 62
rect 7 66 13 70
rect -118 56 -108 60
rect -91 56 -86 64
rect -118 43 -106 56
rect -104 47 -96 56
rect -104 45 -101 47
rect -99 45 -96 47
rect -104 43 -96 45
rect -94 54 -86 56
rect -94 52 -91 54
rect -89 52 -86 54
rect -94 47 -86 52
rect -94 45 -91 47
rect -89 45 -86 47
rect -94 43 -86 45
rect -84 62 -77 64
rect -84 60 -81 62
rect -79 60 -77 62
rect -84 55 -77 60
rect -84 53 -81 55
rect -79 53 -77 55
rect -84 51 -77 53
rect 7 55 12 66
rect -84 43 -79 51
rect 7 43 14 55
rect 16 49 21 55
rect 16 47 23 49
rect 16 45 19 47
rect 21 45 23 47
rect 16 43 23 45
<< alu1 >>
rect -141 72 -73 77
rect -141 70 -110 72
rect -108 70 -102 72
rect -100 70 -73 72
rect -141 69 -73 70
rect 3 72 31 77
rect 3 70 9 72
rect 11 70 19 72
rect 21 70 31 72
rect 3 69 31 70
rect -137 63 -124 64
rect -137 61 -131 63
rect -129 61 -124 63
rect -137 59 -124 61
rect -137 50 -133 59
rect -92 54 -88 56
rect -92 52 -91 54
rect -89 52 -88 54
rect -92 47 -88 52
rect 7 62 19 64
rect 7 60 16 62
rect 18 60 19 62
rect 7 58 19 60
rect 7 57 11 58
rect -36 53 11 57
rect -92 45 -91 47
rect -89 45 -77 47
rect -92 43 -77 45
rect -122 38 -108 39
rect -122 36 -112 38
rect -110 36 -108 38
rect -122 35 -108 36
rect -122 27 -116 35
rect -81 31 -77 43
rect -36 31 -30 53
rect 7 50 11 53
rect 15 47 23 48
rect 15 45 19 47
rect 21 45 23 47
rect 15 44 23 45
rect 15 40 19 44
rect -90 27 -30 31
rect 7 34 19 40
rect 7 29 13 34
rect 7 27 9 29
rect 11 27 13 29
rect -90 23 -86 27
rect 7 26 13 27
rect -100 22 -86 23
rect -100 20 -98 22
rect -96 20 -86 22
rect -100 19 -86 20
rect -141 12 -73 13
rect -141 10 -134 12
rect -132 10 -73 12
rect -141 5 -73 10
rect 3 12 31 13
rect 3 10 10 12
rect 12 10 18 12
rect 20 10 31 12
rect 3 5 31 10
<< ptie >>
rect -136 12 -130 14
rect -136 10 -134 12
rect -132 10 -130 12
rect -136 8 -130 10
rect 8 12 22 17
rect 8 10 10 12
rect 12 10 18 12
rect 20 10 22 12
rect 8 8 22 10
<< ntie >>
rect -112 72 -98 74
rect -112 70 -110 72
rect -108 70 -102 72
rect -100 70 -98 72
rect -112 68 -98 70
rect 17 72 23 74
rect 17 70 19 72
rect 21 70 23 72
rect 17 67 23 70
<< nmos >>
rect -126 24 -124 31
rect 14 25 16 31
rect -113 18 -111 25
rect -103 18 -101 25
rect -93 16 -91 25
rect -86 16 -84 25
<< pmos >>
rect -120 43 -118 64
rect -106 43 -104 56
rect -96 43 -94 56
rect -86 43 -84 64
rect 14 43 16 55
<< polyct0 >>
rect -98 61 -96 63
rect -88 36 -86 38
<< polyct1 >>
rect -131 61 -129 63
rect 16 60 18 62
rect -112 36 -110 38
<< ndifct0 >>
rect -131 27 -129 29
rect 19 27 21 29
rect -120 20 -118 22
rect -108 20 -106 22
rect -81 18 -79 20
<< ndifct1 >>
rect 9 27 11 29
rect -98 20 -96 22
<< ntiect1 >>
rect -110 70 -108 72
rect -102 70 -100 72
rect 19 70 21 72
<< ptiect1 >>
rect -134 10 -132 12
rect 10 10 12 12
rect 18 10 20 12
<< pdifct0 >>
rect -125 45 -123 47
rect -115 60 -113 62
rect -101 45 -99 47
rect -81 60 -79 62
rect -81 53 -79 55
<< pdifct1 >>
rect 9 70 11 72
rect -91 52 -89 54
rect -91 45 -89 47
rect 19 45 21 47
<< alu0 >>
rect -117 62 -111 69
rect -117 60 -115 62
rect -113 60 -111 62
rect -117 59 -111 60
rect -107 63 -78 64
rect -107 61 -98 63
rect -96 62 -78 63
rect -96 61 -81 62
rect -107 60 -81 61
rect -79 60 -78 62
rect -107 55 -103 60
rect -126 51 -103 55
rect -126 47 -122 51
rect -132 45 -125 47
rect -123 45 -122 47
rect -132 43 -122 45
rect -103 47 -97 48
rect -103 45 -101 47
rect -99 45 -97 47
rect -132 29 -128 43
rect -103 39 -97 45
rect -82 55 -78 60
rect -82 53 -81 55
rect -79 53 -78 55
rect -82 51 -78 53
rect -132 27 -131 29
rect -129 27 -128 29
rect -103 38 -84 39
rect -103 36 -88 38
rect -86 36 -84 38
rect -103 35 -84 36
rect -103 31 -99 35
rect -109 27 -99 31
rect -132 25 -128 27
rect -122 22 -116 23
rect -122 20 -120 22
rect -118 20 -116 22
rect -122 13 -116 20
rect -109 22 -105 27
rect 17 29 23 30
rect 17 27 19 29
rect 21 27 23 29
rect -109 20 -108 22
rect -106 20 -105 22
rect -109 18 -105 20
rect -82 20 -78 22
rect -82 18 -81 20
rect -79 18 -78 20
rect -82 13 -78 18
rect 17 13 23 27
<< labels >>
rlabel alu1 9 33 9 33 6 z
rlabel alu1 17 9 17 9 6 vss
rlabel alu1 17 41 17 41 6 z
rlabel alu1 17 73 17 73 6 vdd
rlabel alu0 -124 49 -124 49 6 bn
rlabel alu0 -130 36 -130 36 6 bn
rlabel alu0 -107 24 -107 24 6 an
rlabel alu0 -100 41 -100 41 6 an
rlabel alu0 -94 37 -94 37 6 an
rlabel alu0 -80 57 -80 57 6 bn
rlabel alu0 -93 62 -93 62 6 bn
rlabel alu1 -135 57 -135 57 6 b
rlabel alu1 -127 61 -127 61 6 b
rlabel alu1 -119 33 -119 33 6 a
rlabel polyct1 -111 37 -111 37 6 a
rlabel alu1 -107 9 -107 9 6 vss
rlabel alu1 -107 73 -107 73 6 vdd
<< end >>
