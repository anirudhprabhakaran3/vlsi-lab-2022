magic
tech scmos
timestamp 1663602325
<< polysilicon >>
rect -2 10 0 12
rect -2 1 0 6
rect -5 -1 0 1
rect -2 -6 0 -1
rect -2 -12 0 -10
<< ndiffusion >>
rect -4 -10 -2 -6
rect 0 -10 2 -6
<< pdiffusion >>
rect -4 6 -2 10
rect 0 6 2 10
<< metal1 >>
rect -8 13 6 16
rect -8 10 -5 13
rect 3 -6 6 6
rect -8 -14 -5 -10
rect -8 -17 6 -14
<< ntransistor >>
rect -2 -10 0 -6
<< ptransistor >>
rect -2 6 0 10
<< polycontact >>
rect -9 -2 -5 2
<< ndcontact >>
rect -8 -10 -4 -6
rect 2 -10 6 -6
<< pdcontact >>
rect -8 6 -4 10
rect 2 6 6 10
<< end >>
