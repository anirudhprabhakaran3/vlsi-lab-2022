* NMOS Capacitive Load Inverter

.include ./t14y_tsmc_025_level3.txt

m1 vout vin 0 0 cmosn l=0.5u w=10u
r1 vdd vout 10000
c1 ctop 0 0.1p

v_dd vdd 0 5
v_ctop vout ctop 0
v_in vin 0 PULSE(0 5 0 0.0001n 0.0001n 10m 20m)

.control
        tran 0.001m 100m
        setplot tran1
	plot vin
        plot vout
	plot ctop
        plot -v_dd#branch
	plot -v_ctop#branch
	plot ((1e11*ctop)/(3.14159))
.endc

.end
