* rc simulation




* print output
.op

.control
	
.endc

.end
