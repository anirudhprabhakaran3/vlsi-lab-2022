* nmos characteristics

.include ./t14y_tsmc_025_level3.txt
  
m1 vdd in 0 0 cmosn l=1u w=0.5u 

v_dd vdd 0 3.3 
v_in in 0 3.3 

.control
dc temp -50 125 25
run
setplot dc1
plot (v_in-v_dd)

dc temp -50 125 25
run
setplot dc2
plot (v_in-v_dd)

.end

