magic
tech scmos
timestamp 1666710525
<< pwell >>
rect 0 8 32 32
<< nwell >>
rect 0 32 32 72
<< polysilicon >>
rect 15 50 17 52
rect 15 21 17 38
rect 15 13 17 15
<< ndiffusion >>
rect 0 20 15 21
rect 0 16 5 20
rect 9 16 15 20
rect 0 15 15 16
rect 17 20 32 21
rect 17 16 23 20
rect 27 16 32 20
rect 17 15 32 16
<< pdiffusion >>
rect 0 45 15 50
rect 0 41 5 45
rect 9 41 15 45
rect 0 38 15 41
rect 17 45 32 50
rect 17 41 23 45
rect 27 41 32 45
rect 17 38 32 41
<< metal1 >>
rect 0 64 32 72
rect 5 45 9 64
rect 23 20 27 41
rect 5 8 9 16
rect 0 0 32 8
<< ntransistor >>
rect 15 15 17 21
<< ptransistor >>
rect 15 38 17 50
<< polycontact >>
rect 11 25 15 29
<< ndcontact >>
rect 5 16 9 20
rect 23 16 27 20
<< pdcontact >>
rect 5 41 9 45
rect 23 41 27 45
<< labels >>
rlabel polycontact 13 27 13 27 1 a
rlabel metal1 25 27 25 27 1 output
rlabel metal1 16 4 16 4 1 vss
rlabel metal1 16 68 16 68 5 vdd
<< end >>
