magic
tech scmos
timestamp 1666714927
<< pwell >>
rect 0 29 28 32
rect 0 8 32 29
rect 18 6 32 8
<< nwell >>
rect 0 44 32 64
rect 0 32 28 44
<< polysilicon >>
rect 5 60 7 62
rect 23 60 25 62
rect 5 23 7 44
rect 23 23 25 44
rect 5 12 7 14
rect 23 12 25 14
<< ndiffusion >>
rect 4 14 5 23
rect 7 14 18 23
rect 22 14 23 23
rect 25 14 28 23
<< pdiffusion >>
rect 4 44 5 60
rect 7 54 23 60
rect 7 50 12 54
rect 16 50 23 54
rect 7 44 23 50
rect 25 44 28 60
<< metal1 >>
rect 0 64 32 72
rect 0 60 4 64
rect 28 30 32 44
rect 18 26 32 30
rect 18 23 22 26
rect 0 8 4 14
rect 28 8 32 14
rect 0 0 32 8
<< ntransistor >>
rect 5 14 7 23
rect 23 14 25 23
<< ptransistor >>
rect 5 44 7 60
rect 23 44 25 60
<< polycontact >>
rect 1 37 5 41
rect 19 37 23 41
<< ndcontact >>
rect 0 14 4 23
rect 18 14 22 23
rect 28 14 32 23
<< pdcontact >>
rect 0 44 4 60
rect 28 44 32 60
<< nsubstratencontact >>
rect 12 50 16 54
<< labels >>
rlabel metal1 15 68 15 68 5 vdd
rlabel polycontact 3 39 3 39 3 a
rlabel polycontact 21 39 21 39 1 b
rlabel metal1 15 3 15 3 1 vss
rlabel metal1 30 28 30 28 7 output
rlabel nsubstratencontact 14 52 14 52 1 psub
<< end >>
