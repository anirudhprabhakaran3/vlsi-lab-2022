* nmos characteristics

* include the model files
.include ./t14y_tsmc_025_level3.txt
  
* netlist
* m_instance_name drain_node gate_node source_node bulk_substrate_node model_name L=length W=width

m1 vdd in 0 0 cmosn w=1u 

v_dd vdd 0 3.3 
v_in in 0 3.3 

.control
        let nmoslength = 0.5u
        let plotnum = 1
        dowhile nmoslength <= 10u

                alter @m1[l] = nmoslength
	
                dc v_in 0 3.3 0.1 v_dd 0 3.3 1
                run
                setplot dc$plotnum
                plot -v_dd#branch

                let plotnum = plotnum + 1
                let nmoslength = nmoslength + 1u
        end
.endc

.end

