* SPICE3 file created from new_invertor.ext - technology: scmos

.include ./t14y_tsmc_025_level3.txt

.option scale=1u

M1000 out in vdd vdd cmosp w=8 l=2
+  ad=40 pd=26 as=40 ps=26
M1001 out in vss Gnd cmosn w=4 l=2
+  ad=20 pd=18 as=20 ps=18
* C0 vss Gnd 2.26fF
* C1 in Gnd 4.68fF


v_dd vdd Gnd 5
v_in in Gnd PULSE(0 5 0 0 2 10 20)
v_gnd Gnd 0 20

.control
	tran 0.1 40
	setplot tran1
	plot in out
.endc

.end
