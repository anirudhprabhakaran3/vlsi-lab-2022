magic
tech scmos
timestamp 1666020471
<< ab >>
rect -87 5 -23 77
rect 5 5 29 77
<< nwell >>
rect -11 82 -10 97
rect -92 37 34 82
<< pwell >>
rect -92 0 34 37
<< poly >>
rect -77 67 -66 69
rect -77 65 -75 67
rect -81 63 -75 65
rect -68 64 -66 67
rect -81 61 -79 63
rect -77 61 -75 63
rect -81 59 -75 61
rect -48 63 -42 65
rect -34 64 -32 69
rect -48 61 -46 63
rect -44 61 -42 63
rect -54 56 -52 61
rect -48 59 -42 61
rect -44 56 -42 59
rect 14 62 20 64
rect 14 60 16 62
rect 18 60 20 62
rect 14 58 20 60
rect 14 55 16 58
rect -68 40 -66 43
rect -54 40 -52 43
rect -74 38 -66 40
rect -62 38 -52 40
rect -74 31 -72 38
rect -62 36 -60 38
rect -58 36 -56 38
rect -62 34 -56 36
rect -61 25 -59 34
rect -44 30 -42 43
rect -34 40 -32 43
rect -38 38 -32 40
rect -38 36 -36 38
rect -34 36 -32 38
rect -38 34 -32 36
rect -51 25 -49 30
rect -44 28 -39 30
rect -41 25 -39 28
rect -34 25 -32 34
rect 14 31 16 43
rect -74 10 -72 24
rect -61 14 -59 18
rect -51 10 -49 18
rect 14 20 16 25
rect -41 11 -39 16
rect -34 11 -32 16
rect -74 8 -49 10
<< ndif >>
rect -81 29 -74 31
rect -81 27 -79 29
rect -77 27 -74 29
rect -81 24 -74 27
rect -72 25 -63 31
rect 7 29 14 31
rect 7 27 9 29
rect 11 27 14 29
rect 7 25 14 27
rect 16 29 23 31
rect 16 27 19 29
rect 21 27 23 29
rect 16 25 23 27
rect -72 24 -61 25
rect -70 22 -61 24
rect -70 20 -68 22
rect -66 20 -61 22
rect -70 18 -61 20
rect -59 22 -51 25
rect -59 20 -56 22
rect -54 20 -51 22
rect -59 18 -51 20
rect -49 22 -41 25
rect -49 20 -46 22
rect -44 20 -41 22
rect -49 18 -41 20
rect -46 16 -41 18
rect -39 16 -34 25
rect -32 20 -25 25
rect -32 18 -29 20
rect -27 18 -25 20
rect -32 16 -25 18
<< pdif >>
rect 7 72 13 74
rect 7 70 9 72
rect 11 70 13 72
rect -73 49 -68 64
rect -75 47 -68 49
rect -75 45 -73 47
rect -71 45 -68 47
rect -75 43 -68 45
rect -66 62 -56 64
rect -66 60 -63 62
rect -61 60 -56 62
rect 7 66 13 70
rect -66 56 -56 60
rect -39 56 -34 64
rect -66 43 -54 56
rect -52 47 -44 56
rect -52 45 -49 47
rect -47 45 -44 47
rect -52 43 -44 45
rect -42 54 -34 56
rect -42 52 -39 54
rect -37 52 -34 54
rect -42 47 -34 52
rect -42 45 -39 47
rect -37 45 -34 47
rect -42 43 -34 45
rect -32 62 -25 64
rect -32 60 -29 62
rect -27 60 -25 62
rect -32 55 -25 60
rect -32 53 -29 55
rect -27 53 -25 55
rect -32 51 -25 53
rect 7 55 12 66
rect -32 43 -27 51
rect 7 43 14 55
rect 16 49 21 55
rect 16 47 23 49
rect 16 45 19 47
rect 21 45 23 47
rect 16 43 23 45
<< alu1 >>
rect -89 72 -21 77
rect -89 70 -58 72
rect -56 70 -50 72
rect -48 70 -21 72
rect -89 69 -21 70
rect 3 72 31 77
rect 3 70 9 72
rect 11 70 19 72
rect 21 70 31 72
rect 3 69 31 70
rect -85 63 -72 64
rect -85 61 -79 63
rect -77 61 -72 63
rect -85 59 -72 61
rect -85 50 -81 59
rect -40 54 -36 56
rect -40 52 -39 54
rect -37 52 -36 54
rect -40 47 -36 52
rect -11 62 19 64
rect -11 60 16 62
rect 18 60 19 62
rect -40 45 -39 47
rect -37 45 -25 47
rect -40 43 -25 45
rect -70 38 -56 39
rect -70 36 -60 38
rect -58 36 -56 38
rect -70 35 -56 36
rect -70 27 -64 35
rect -29 31 -25 43
rect -11 31 -7 60
rect 7 58 19 60
rect 7 50 11 58
rect 15 47 23 48
rect 15 45 19 47
rect 21 45 23 47
rect 15 44 23 45
rect 15 40 19 44
rect -38 27 -7 31
rect 7 34 19 40
rect 7 29 13 34
rect 7 27 9 29
rect 11 27 13 29
rect -38 23 -34 27
rect 7 26 13 27
rect -48 22 -34 23
rect -48 20 -46 22
rect -44 20 -34 22
rect -48 19 -34 20
rect -89 12 -21 13
rect -89 10 -82 12
rect -80 10 -21 12
rect -89 5 -21 10
rect 3 12 31 13
rect 3 10 10 12
rect 12 10 18 12
rect 20 10 31 12
rect 3 5 31 10
<< ptie >>
rect -84 12 -78 14
rect -84 10 -82 12
rect -80 10 -78 12
rect -84 8 -78 10
rect 8 12 22 17
rect 8 10 10 12
rect 12 10 18 12
rect 20 10 22 12
rect 8 8 22 10
<< ntie >>
rect -60 72 -46 74
rect -60 70 -58 72
rect -56 70 -50 72
rect -48 70 -46 72
rect -60 68 -46 70
rect 17 72 23 74
rect 17 70 19 72
rect 21 70 23 72
rect 17 67 23 70
<< nmos >>
rect -74 24 -72 31
rect 14 25 16 31
rect -61 18 -59 25
rect -51 18 -49 25
rect -41 16 -39 25
rect -34 16 -32 25
<< pmos >>
rect -68 43 -66 64
rect -54 43 -52 56
rect -44 43 -42 56
rect -34 43 -32 64
rect 14 43 16 55
<< polyct0 >>
rect -46 61 -44 63
rect -36 36 -34 38
<< polyct1 >>
rect -79 61 -77 63
rect 16 60 18 62
rect -60 36 -58 38
<< ndifct0 >>
rect -79 27 -77 29
rect 19 27 21 29
rect -68 20 -66 22
rect -56 20 -54 22
rect -29 18 -27 20
<< ndifct1 >>
rect 9 27 11 29
rect -46 20 -44 22
<< ntiect1 >>
rect -58 70 -56 72
rect -50 70 -48 72
rect 19 70 21 72
<< ptiect1 >>
rect -82 10 -80 12
rect 10 10 12 12
rect 18 10 20 12
<< pdifct0 >>
rect -73 45 -71 47
rect -63 60 -61 62
rect -49 45 -47 47
rect -29 60 -27 62
rect -29 53 -27 55
<< pdifct1 >>
rect 9 70 11 72
rect -39 52 -37 54
rect -39 45 -37 47
rect 19 45 21 47
<< alu0 >>
rect -65 62 -59 69
rect -65 60 -63 62
rect -61 60 -59 62
rect -65 59 -59 60
rect -55 63 -26 64
rect -55 61 -46 63
rect -44 62 -26 63
rect -44 61 -29 62
rect -55 60 -29 61
rect -27 60 -26 62
rect -55 55 -51 60
rect -74 51 -51 55
rect -74 47 -70 51
rect -80 45 -73 47
rect -71 45 -70 47
rect -80 43 -70 45
rect -51 47 -45 48
rect -51 45 -49 47
rect -47 45 -45 47
rect -80 29 -76 43
rect -51 39 -45 45
rect -30 55 -26 60
rect -30 53 -29 55
rect -27 53 -26 55
rect -30 51 -26 53
rect -80 27 -79 29
rect -77 27 -76 29
rect -51 38 -32 39
rect -51 36 -36 38
rect -34 36 -32 38
rect -51 35 -32 36
rect -51 31 -47 35
rect -57 27 -47 31
rect -80 25 -76 27
rect -70 22 -64 23
rect -70 20 -68 22
rect -66 20 -64 22
rect -70 13 -64 20
rect -57 22 -53 27
rect 17 29 23 30
rect 17 27 19 29
rect 21 27 23 29
rect -57 20 -56 22
rect -54 20 -53 22
rect -57 18 -53 20
rect -30 20 -26 22
rect -30 18 -29 20
rect -27 18 -26 20
rect -30 13 -26 18
rect 17 13 23 27
<< labels >>
rlabel alu1 9 33 9 33 6 z
rlabel alu1 17 9 17 9 6 vss
rlabel alu1 17 41 17 41 6 z
rlabel alu1 17 73 17 73 6 vdd
rlabel alu0 -72 49 -72 49 6 bn
rlabel alu0 -78 36 -78 36 6 bn
rlabel alu0 -55 24 -55 24 6 an
rlabel alu0 -48 41 -48 41 6 an
rlabel alu0 -42 37 -42 37 6 an
rlabel alu0 -28 57 -28 57 6 bn
rlabel alu0 -41 62 -41 62 6 bn
rlabel alu1 -83 57 -83 57 6 b
rlabel alu1 -75 61 -75 61 6 b
rlabel alu1 -67 33 -67 33 6 a
rlabel polyct1 -59 37 -59 37 6 a
rlabel alu1 -55 9 -55 9 6 vss
rlabel alu1 -55 73 -55 73 6 vdd
<< end >>
