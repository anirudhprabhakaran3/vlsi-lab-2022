* nmos characteristics

.include ./t14y_tsmc_025_level3.txt
  
m1 vdd in 1 0 cmosn l=1u w=0.5u
m2 vdd2 in2 5 0 cmosn l=1u w=0.5u  

v_dd vdd 0 3.3 
v_in in 0 3.3 

v_dd2 vdd2 0 3.3
v_in2 in2 0 3.3

.control
dc v_in 0 3.3 0.1 v_dd 0 3.3 1
run
setplot dc1
plot -v_dd#branch

dc v_dd 0 3.3 .1 v_in 0 3.3  .1
run
setplot dc2
plot -v_dd#branch

dc v_in2 0 3.3 0.1 v_dd2 0 3.3 1
run
setplot dc3
plot -v_dd2#branch

dc v_dd2 0 3.3 0.1 v_in2 0 3.3 1
run
setplot dc4
plot -v_dd2#branch
.endc

.end

