magic
tech scmos
timestamp 1199202227
<< ab >>
rect 0 0 24 72
<< nwell >>
rect -5 32 29 77
<< pwell >>
rect -5 -5 29 32
<< poly >>
rect 9 57 15 59
rect 9 55 11 57
rect 13 55 15 57
rect 9 53 15 55
rect 9 50 11 53
rect 9 26 11 38
rect 9 15 11 20
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 20 9 22
rect 11 24 18 26
rect 11 22 14 24
rect 16 22 18 24
rect 11 20 18 22
<< pdif >>
rect 2 67 8 69
rect 2 65 4 67
rect 6 65 8 67
rect 2 61 8 65
rect 2 50 7 61
rect 2 38 9 50
rect 11 44 16 50
rect 11 42 18 44
rect 11 40 14 42
rect 16 40 18 42
rect 11 38 18 40
<< alu1 >>
rect -2 67 26 72
rect -2 65 4 67
rect 6 65 14 67
rect 16 65 26 67
rect -2 64 26 65
rect 2 57 14 59
rect 2 55 11 57
rect 13 55 14 57
rect 2 53 14 55
rect 2 45 6 53
rect 10 42 18 43
rect 10 40 14 42
rect 16 40 18 42
rect 10 39 18 40
rect 10 35 14 39
rect 2 29 14 35
rect 2 24 8 29
rect 2 22 4 24
rect 6 22 8 24
rect 2 21 8 22
rect -2 7 26 8
rect -2 5 5 7
rect 7 5 13 7
rect 15 5 26 7
rect -2 0 26 5
<< ptie >>
rect 3 7 17 12
rect 3 5 5 7
rect 7 5 13 7
rect 15 5 17 7
rect 3 3 17 5
<< ntie >>
rect 12 67 18 69
rect 12 65 14 67
rect 16 65 18 67
rect 12 62 18 65
<< nmos >>
rect 9 20 11 26
<< pmos >>
rect 9 38 11 50
<< polyct1 >>
rect 11 55 13 57
<< ndifct0 >>
rect 14 22 16 24
<< ndifct1 >>
rect 4 22 6 24
<< ntiect1 >>
rect 14 65 16 67
<< ptiect1 >>
rect 5 5 7 7
rect 13 5 15 7
<< pdifct1 >>
rect 4 65 6 67
rect 14 40 16 42
<< alu0 >>
rect 12 24 18 25
rect 12 22 14 24
rect 16 22 18 24
rect 12 8 18 22
<< labels >>
rlabel alu1 4 28 4 28 6 z
rlabel alu1 4 52 4 52 6 a
rlabel alu1 12 4 12 4 6 vss
rlabel alu1 12 36 12 36 6 z
rlabel alu1 12 68 12 68 6 vdd
rlabel polyct1 12 56 12 56 6 a
<< end >>
